package constant;
	parameter INST_SIZE = 15;
	parameter BRAM_SIZE = 19;
endpackage
